`ifndef PARAM_SVH
`define PARAM_SVH

`define BIT_WIDTH 32

`endif  // PARAM_SVH
